LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY PC IS
	PORT(
		CLK :							IN		STD_LOGIC;
		RESET :						IN		STD_LOGIC;
		IN_PC :						IN 	STD_LOGIC_VECTOR(31 DOWNTO 0);
		OUT_PC :						OUT	STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END PC;

ARCHITECTURE ARC_PC OF PC IS
	
BEGIN
	PROCESS(CLK, RESET)
	BEGIN
		IF RESET = '1' THEN
			OUT_A <= X"00400000";								--Para utilizar com o MARS
		ELSIF	CLK'EVENT AND CLK = '1' THEN
			OUT_A <= IN_A;
		END IF;
	END PROCESS;
END ARC_PC;